module dist_mem_gen_0 (input [11:0] a,
                       input [15:0] d,
                       input clk,
                       we,
                       output [15:0] spo);

endmodule
