module alu #(parameter WIDTH = 32)
    (input [WIDTH - 1: 0] a,
     input [WIDTH - 1: 0] b,      // 两操作数
     input [2:0] s,               // 功能选择
     output reg [WIDTH - 1: 0] y, // 运算结果
     output reg [2:0] f);         // 标志

    wire a_s, b_s;
    assign a_s = ~a[WIDTH - 1];
    assign b_s = ~b[WIDTH - 1];

    always @(*) begin
        f = 3'b000;
        y = 0;
        case (s)
            3'b000:
                y = a - b;
            3'b001:
                y = a + b;
            3'b010:
                y = a & b;
            3'b011:
                y = a | b;
            3'b100:
                y = a ^ b;
            3'b101:
                y = a >> b;
            3'b110:
                y = a << b;
            3'b111:
                y = ($signed(a)) >>> b;       // signed
        endcase
        if (s == 3'b000) begin
            f[0] = (y == 0 ? 1'b1 :1'b0);
            f[1] = {a_s, a} < {b_s, b} ? 1'b1 : 1'b0;
            f[2] = (a < b ? 1'b1 :1'b0);
        end
    end
endmodule
